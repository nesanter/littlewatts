Punk v2 (Class-A Amplifier)
****
* Author: Noah Santer (santerkrupp@gmail.com)
****

*** Parameters ***
.param rail_voltage = 24V
.param input_voltage = 400mV
.param input_frequency = 1KHz

.param Rq = 1Kohm
.param Rg = 2.2Kohm

*** Supply ***
Bvcc vcc 0 V = rail_voltage
.save @bvcc[i]

*** Signal ***
Vsig sig 0 dc 0V ac 1V sine(0V input_voltage input_frequency)
.save v(sig)

*** Load ***
Rload output 0 8ohm
.save v(output)
.save @rload[p]

*** Input ***
R1 sig 100 6.8Kohm
R2 100 vcc 10Kohm

Q1 101 100 102 Q2N3904
Q2 103 nfb 104 Q2N3904

Q3 101 103 vcc Q2N3906
Q4 103 103 vcc Q2N3906

R3 102 105 0ohm
R4 104 105 0ohm


Q5 105 106 107 Q2N2222A
Q6 106 107 0 Q2N2222A
R5 106 vcc 220Kohm
R6 107 0 100ohm

*** VAS ***
Q7 0 101 108 Q2N3906
R7 108 vcc 1Kohm
Q8 109 108 vcc Q2N3906
Q9 109 106 110 Q2N3904
R8 110 0 100ohm
C1 101 109 10pF

*** Drive ***
R9 vcc h 0ohm
R10 l 0 0.0ohm
Q10a h 109 112ha QC4883A
Q10b h 109 112hb QC4883A
Q10c h 109 112hc QC4883A
*Q10d h 109 112hd QC4883A
Rswamp1 112ha 112 0.22ohm
Rswamp2 112hb 112 0.22ohm
Rswamp3 112hc 112 0.22ohm
*Rswamp4 112hd 112 0.22ohm

Q11a 112 113 la QC4883A
Q11b 112 113 lb QC4883A
Q11c 112 113 lc QC4883A
*Q11d 112 113 ld QC4883A
Rswamp5 la l 0.22ohm
Rswamp6 lb l 0.22ohm
Rswamp7 lc l 0.22ohm
*Rswamp8 ld l 0.22ohm

C2 h 113 100pF
R11 vcc 115 100ohm
R12 115b 0 330ohm
R13 113b 113 Rq
Q12 115 113b 115b Q2N3906

.save @q10a[p]
.save @q11a[p]

*** Ouput & NFB ***
R14 112 nfb 100Kohm
R15 nfb 116 Rg
C3 116 0 220uF

C4 112 output 2200uF

*** Analysis ***
.control
tran 10u 1

fourier 1K v(output)

meas tran rmspout rms @rload[p]
meas tran rmsivcc rms @bvcc[i]
meas tran avgpq10a avg @q10a[p]
meas tran avgpq11 avg @q11a[p]
.endc

*** Models ***
.MODEL Q2N2222A npn (
+IS=3.88184e-14 BF=929.846 NF=1.10496 VAF=16.5003
+IKF=0.019539 ISE=1.0168e-11 NE=1.94752 BR=48.4545
+NR=1.07004 VAR=40.538 IKR=0.19539 ISC=1.0168e-11
+NC=4 RB=0.1 IRB=0.1 RBM=0.1
+RE=0.0001 RC=0.426673 XTB=0.1 XTI=1
+EG=1.05 CJE=2.23677e-11 VJE=0.582701 MJE=0.63466
+TF=4.06711e-10 XTF=3.92912 VTF=17712.6 ITF=0.4334
+CJC=2.23943e-11 VJC=0.576146 MJC=0.632796 XCJC=1
+FC=0.170253 CJS=0 VJS=0.75 MJS=0.5
+TR=1e-07 PTF=0 KF=0 AF=1 )

.MODEL QMJL3281A npn IS=9.8145e-12 BF=438.0 NF=1.00 VAF=38 IKF=19.0 ISE=1.0e-12 NE=1.1237388682 BR=4.98985 NR=1.09511 VAR=4.32026 IKR=4.37516 ISC=3.25e-13 NC=3.96875 RB=3.997 RE=0.00 RC=0.06 XTB=0.115253 XTI=1.03146 EG=1.11986 CJE=1.144e-08 VJE=0.468574 MJE=0.34957 TF=2.6769e-9 XTF=7500 VTF=3.0 ITF=1000 CJC=1.093685e-9 VJC=0.623643 MJC=0.482111 XCJC=0.959922 FC=0.1 CJS=0 VJS=0.75 MJS=0.5 TR=1e-07 PTF=0 KF=0 AF=1 Vceo=200

.model QC4883A NPN (level=2 Bf=140 Ikf=100 Is=600f Vaf=100 
+ Rb=1.7 Re=105m RC=0 Isc=150f
+ Cje=1.2n Cjc=72p Tf=875p Vtf=1.2 Itf=1
+ Br=2 Var=22.9 Ikr=36 TR=85n
+ Xtb=0.34 Xtf=1.36 )

.MODEL Q2N3904 npn IS=3.5e-15 BF=160 VAF=400 IKF=0.15 ISE=4e-16 NE=1.26 NF=1 RB=30.1 RC=1 RE=0.1 CJE=15e-12 MJE=0.25 VJE=0.75 CJC=3.6e-12 MJC=0.30 VJC=0.75 FC=0.5 TF=380e-12 XTF=30 VTF=4 ITF=0.4 TR=240e-9 BR=0.7 IKR=0 EG=1.1 XTB=1.5 XTI=3 NC=2 ISC=0
.MODEL Q2N3906 pnp IS=10e-15 BF=180 VAF=40 IKF=0.6 ISE=30e-15 NE=1.5 NF=1 RB=33 RC=1 RE=0.1 CJE=12e-12 MJE=0.7 VJE=1.0 CJC=12e-12 MJC=0.7 VJC=1.0 FC=0.5 TF=550e-12 XTF=20000 VTF=10 ITF=3.5 TR=10e-9 BR=4 IKR=11 EG=1.1 XTB=1.5 XTI=3 NC=15.5 ISC=0.5e-15 VAR=100 NK=1.0

.MODEL QA1859A pnp (Bf=162 IKF=10 Is=500f Vaf=300 
+ Rb=0 Re=0 Rc=90m Rco=3.25 Ibc=150f Vo=120 Gamma=22n
+ Cje=1.5n Cjc=72p Tf=1.9n Vtf=1.9 Itf=1 Qco=8p
+ Br=2 Ikr=10 Var=23 Tr=188.8n
+ Xtb=0.138 Xtf=5)

.end
